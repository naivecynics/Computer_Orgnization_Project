module cpu_top(
    input fpga_rst,     // active high
    input fpga_clk,

    input start_pg,
    input rx,
    output tx
);



endmodule