`timescale 1ns / 1ps

module instr_decoder(   
    input [31:0] instr;
    output [6:0] opcode;
    