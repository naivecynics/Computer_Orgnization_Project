`timescale 1ns/1ps

module debounce(
    input clk,
    input rst_n;
    input key_in,
    output key_out
);


endmodule